module processor;


endmodule 
